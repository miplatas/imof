library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Inversor is

generic(
    delay: integer := 15 -- max delay 19 pulsos
    );


    Port ( clk         : in  STD_LOGIC;
           start      : in STD_LOGIC;
           reset, mode      : in STD_LOGIC;
           freq_carrier  : in  STD_LOGIC_VECTOR(15 downto 0); 
           freq_sine  : in  STD_LOGIC_VECTOR(15 downto 0); 
           LED    : out STD_LOGIC_VECTOR(15 downto 0);
           igbt    : out STD_LOGIC_VECTOR(5 downto 0);
           enable : out std_logic
           ); 
end Inversor;

architecture Behavioral of Inversor is

signal state_reg, state_next, enable_reg, enable_next : std_logic;

type sine_table_type is array(0 to 4095) of unsigned(11 downto 0); -- 12 bits de resolución
constant sine_table: sine_table_type := (    
"011111111111", "011111111100", "011111111001", "011111110110", "011111110011", "011111110000", "011111101101", "011111101010", "011111100111", "011111100100", "011111100000", "011111011101", "011111011010", "011111010111", "011111010100", "011111010001", "011111001110", "011111001011", "011111001000", "011111000100", "011111000001", "011110111110", "011110111011", "011110111000", "011110110101", "011110110010", "011110101111", "011110101100", "011110101000", "011110100101", "011110100010", "011110011111", "011110011100", "011110011001", "011110010110", "011110010011", "011110010000", "011110001100", "011110001001", "011110000110", "011110000011", "011110000000", "011101111101", "011101111010", "011101110111", "011101110100", "011101110001", "011101101101", "011101101010", "011101100111", "011101100100", "011101100001", "011101011110", "011101011011", "011101011000", "011101010101", "011101010010", "011101001110", "011101001011", "011101001000", "011101000101", "011101000010", "011100111111", "011100111100", "011100111001", "011100110110", "011100110011", "011100101111", "011100101100", "011100101001", "011100100110", "011100100011", "011100100000", "011100011101", "011100011010", "011100010111", "011100010100", "011100010001", "011100001101", "011100001010", "011100000111", "011100000100", "011100000001", "011011111110", "011011111011", "011011111000", "011011110101", "011011110010", "011011101111", "011011101100", "011011101000", "011011100101", "011011100010", "011011011111", "011011011100", "011011011001", "011011010110", "011011010011", "011011010000", "011011001101", "011011001010", "011011000111", "011011000100", "011011000000", "011010111101", "011010111010", "011010110111", "011010110100", "011010110001", "011010101110", "011010101011", "011010101000", "011010100101", "011010100010", "011010011111", "011010011100", "011010011001", "011010010110", "011010010011", "011010001111", "011010001100", "011010001001", "011010000110", "011010000011", "011010000000", "011001111101", "011001111010", "011001110111", "011001110100", "011001110001", "011001101110", "011001101011", "011001101000", "011001100101", "011001100010", "011001011111", "011001011100", "011001011001", "011001010101", "011001010010", "011001001111", "011001001100", "011001001001", "011001000110", "011001000011", "011001000000", "011000111101", "011000111010", "011000110111", "011000110100", "011000110001", "011000101110", "011000101011", "011000101000", "011000100101", "011000100010", "011000011111", "011000011100", "011000011001", "011000010110", "011000010011", "011000010000", "011000001101", "011000001010", "011000000111", "011000000100", "011000000001", "010111111110", "010111111011", "010111111000", "010111110101", "010111110010", "010111101111", "010111101100", "010111101001", "010111100110", "010111100011", "010111100000", "010111011101", "010111011010", "010111010111", "010111010100", "010111010001", "010111001110", "010111001011", "010111001000", "010111000101", "010111000010", "010110111111", "010110111100", "010110111001", "010110110110", "010110110011", "010110110000", "010110101101", "010110101010", "010110100111", "010110100100", "010110100001", "010110011110", "010110011011", "010110011000", "010110010101", "010110010010", "010110001111", "010110001100", "010110001001", "010110000110", "010110000100", "010110000001", "010101111110", "010101111011", "010101111000", "010101110101", "010101110010", "010101101111", "010101101100", "010101101001", "010101100110", "010101100011", "010101100000", "010101011101", "010101011010", "010101010111", "010101010100", "010101010010", "010101001111", "010101001100", "010101001001", "010101000110", "010101000011", "010101000000", "010100111101", "010100111010", "010100110111", "010100110100", "010100110001", "010100101111", "010100101100", "010100101001", "010100100110", "010100100011", "010100100000", "010100011101", "010100011010", "010100010111", "010100010100", "010100010010", "010100001111", "010100001100", "010100001001", "010100000110", "010100000011", "010100000000", "010011111101", "010011111010", "010011111000", "010011110101", "010011110010", "010011101111", "010011101100", "010011101001", "010011100110", "010011100100", "010011100001", "010011011110", "010011011011", "010011011000", "010011010101", "010011010010", "010011010000", "010011001101", "010011001010", "010011000111", "010011000100", "010011000001", "010010111111", "010010111100", "010010111001", "010010110110", "010010110011", "010010110000", "010010101110", "010010101011", "010010101000", "010010100101", "010010100010", "010010011111", "010010011101", "010010011010", "010010010111", "010010010100", "010010010001", "010010001111", "010010001100", "010010001001", "010010000110", "010010000011", "010010000001", "010001111110", "010001111011", "010001111000", "010001110101", "010001110011", "010001110000", "010001101101", "010001101010", "010001101000", "010001100101", "010001100010", "010001011111", "010001011101", "010001011010", "010001010111", "010001010100", "010001010001", "010001001111", "010001001100", "010001001001", "010001000110", "010001000100", "010001000001", "010000111110", "010000111100", "010000111001", "010000110110", "010000110011", "010000110001", "010000101110", "010000101011", "010000101000", "010000100110", "010000100011", "010000100000", "010000011110", "010000011011", "010000011000", "010000010101", "010000010011", "010000010000", "010000001101", "010000001011", "010000001000", "010000000101", "010000000011", "010000000000", "001111111101", "001111111011", "001111111000", "001111110101", "001111110011", "001111110000", "001111101101", "001111101011", "001111101000", "001111100101", "001111100011", "001111100000", "001111011101", "001111011011", "001111011000", "001111010101", "001111010011", "001111010000", "001111001101", "001111001011", "001111001000", "001111000101", "001111000011", "001111000000", "001110111110", "001110111011", "001110111000", "001110110110", "001110110011", "001110110000", "001110101110", "001110101011", "001110101001", "001110100110", "001110100011", "001110100001", "001110011110", "001110011100", "001110011001", "001110010111", "001110010100", "001110010001", "001110001111", "001110001100", "001110001010", "001110000111", "001110000101", "001110000010", "001101111111", "001101111101", "001101111010", "001101111000", "001101110101", "001101110011", "001101110000", "001101101110", "001101101011", "001101101000", "001101100110", "001101100011", "001101100001", "001101011110", "001101011100", "001101011001", "001101010111", "001101010100", "001101010010", "001101001111", "001101001101", "001101001010", "001101001000", "001101000101", "001101000011", "001101000000", "001100111110", "001100111011", "001100111001", "001100110110", "001100110100", "001100110001", "001100101111", "001100101100", "001100101010", "001100101000", "001100100101", "001100100011", "001100100000", "001100011110", "001100011011", "001100011001", "001100010110", "001100010100", "001100010001", "001100001111", "001100001101", "001100001010", "001100001000", "001100000101", "001100000011", "001100000001", "001011111110", "001011111100", "001011111001", "001011110111", "001011110101", "001011110010", "001011110000", "001011101101", "001011101011", "001011101001", "001011100110", "001011100100", "001011100001", "001011011111", "001011011101", "001011011010", "001011011000", "001011010110", "001011010011", "001011010001", "001011001111", "001011001100", "001011001010", "001011001000", "001011000101", "001011000011", "001011000000", "001010111110", "001010111100", "001010111010", "001010110111", "001010110101", "001010110011", "001010110000", "001010101110", "001010101100", "001010101001", "001010100111", "001010100101", "001010100010", "001010100000", "001010011110", "001010011100", "001010011001", "001010010111", "001010010101", "001010010011", "001010010000", "001010001110", "001010001100", "001010001010", "001010000111", "001010000101", "001010000011", "001010000001", "001001111110", "001001111100", "001001111010", "001001111000", "001001110101", "001001110011", "001001110001", "001001101111", "001001101101", "001001101010", "001001101000", "001001100110", "001001100100", "001001100010", "001001011111", "001001011101", "001001011011", "001001011001", "001001010111", "001001010100", "001001010010", "001001010000", "001001001110", "001001001100", "001001001010", "001001000111", "001001000101", "001001000011", "001001000001", "001000111111", "001000111101", "001000111011", "001000111000", "001000110110", "001000110100", "001000110010", "001000110000", "001000101110", "001000101100", "001000101010", "001000101000", "001000100101", "001000100011", "001000100001", "001000011111", "001000011101", "001000011011", "001000011001", "001000010111", "001000010101", "001000010011", "001000010001", "001000001111", "001000001101", "001000001011", "001000001000", "001000000110", "001000000100", "001000000010", "001000000000", "000111111110", "000111111100", "000111111010", "000111111000", "000111110110", "000111110100", "000111110010", "000111110000", "000111101110", "000111101100", "000111101010", "000111101000", "000111100110", "000111100100", "000111100010", "000111100000", "000111011110", "000111011100", "000111011010", "000111011000", "000111010110", "000111010101", "000111010011", "000111010001", "000111001111", "000111001101", "000111001011", "000111001001", "000111000111", "000111000101", "000111000011", "000111000001", "000110111111", "000110111101", "000110111100", "000110111010", "000110111000", "000110110110", "000110110100", "000110110010", "000110110000", "000110101110", "000110101100", "000110101011", "000110101001", "000110100111", "000110100101", "000110100011", "000110100001", "000110011111", "000110011110", "000110011100", "000110011010", "000110011000", "000110010110", "000110010100", "000110010011", "000110010001", "000110001111", "000110001101", "000110001011", "000110001010", "000110001000", "000110000110", "000110000100", "000110000010", "000110000001", "000101111111", "000101111101", "000101111011", "000101111010", "000101111000", "000101110110", "000101110100", "000101110011", "000101110001", "000101101111", "000101101101", "000101101100", "000101101010", "000101101000", "000101100110", "000101100101", "000101100011", "000101100001", "000101100000", "000101011110", "000101011100", "000101011010", "000101011001", "000101010111", "000101010101", "000101010100", "000101010010", "000101010000", "000101001111", "000101001101", "000101001011", "000101001010", "000101001000", "000101000110", "000101000101", "000101000011", "000101000010", "000101000000", "000100111110", "000100111101", "000100111011", "000100111001", "000100111000", "000100110110", "000100110101", "000100110011", "000100110001", "000100110000", "000100101110", "000100101101", "000100101011", "000100101010", "000100101000", "000100100110", "000100100101", "000100100011", "000100100010", "000100100000", "000100011111", "000100011101", "000100011100", "000100011010", "000100011000", "000100010111", "000100010101", "000100010100", "000100010010", "000100010001", "000100001111", "000100001110", "000100001100", "000100001011", "000100001001", "000100001000", "000100000111", "000100000101", "000100000100", "000100000010", "000100000001", "000011111111", "000011111110", "000011111100", "000011111011", "000011111001", "000011111000", "000011110111", "000011110101", "000011110100", "000011110010", "000011110001", "000011101111", "000011101110", "000011101101", "000011101011", "000011101010", "000011101000", "000011100111", "000011100110", "000011100100", "000011100011", "000011100010", "000011100000", "000011011111", "000011011110", "000011011100", "000011011011", "000011011010", "000011011000", "000011010111", "000011010110", "000011010100", "000011010011", "000011010010", "000011010000", "000011001111", "000011001110", "000011001100", "000011001011", "000011001010", "000011001000", "000011000111", "000011000110", "000011000101", "000011000011", "000011000010", "000011000001", "000011000000", "000010111110", "000010111101", "000010111100", "000010111011", "000010111001", "000010111000", "000010110111", "000010110110", "000010110101", "000010110011", "000010110010", "000010110001", "000010110000", "000010101111", "000010101101", "000010101100", "000010101011", "000010101010", "000010101001", "000010100111", "000010100110", "000010100101", "000010100100", "000010100011", "000010100010", "000010100001", "000010011111", "000010011110", "000010011101", "000010011100", "000010011011", "000010011010", "000010011001", "000010011000", "000010010111", "000010010101", "000010010100", "000010010011", "000010010010", "000010010001", "000010010000", "000010001111", "000010001110", "000010001101", "000010001100", "000010001011", "000010001010", "000010001001", "000010001000", "000010000111", "000010000110", "000010000101", "000010000100", "000010000011", "000010000010", "000010000001", "000010000000", "000001111111", "000001111110", "000001111101", "000001111100", "000001111011", "000001111010", "000001111001", "000001111000", "000001110111", "000001110110", "000001110101", "000001110100", "000001110011", "000001110010", "000001110001", "000001110000", "000001101111", "000001101110", "000001101101", "000001101100", "000001101100", "000001101011", "000001101010", "000001101001", "000001101000", "000001100111", "000001100110", "000001100101", "000001100101", "000001100100", "000001100011", "000001100010", "000001100001", "000001100000", "000001011111", "000001011111", "000001011110", "000001011101", "000001011100", "000001011011", "000001011010", "000001011010", "000001011001", "000001011000", "000001010111", "000001010110", "000001010110", "000001010101", "000001010100", "000001010011", "000001010011", "000001010010", "000001010001", "000001010000", "000001010000", "000001001111", "000001001110", "000001001101", "000001001101", "000001001100", "000001001011", "000001001010", "000001001010", "000001001001", "000001001000", "000001001000", "000001000111", "000001000110", "000001000110", "000001000101", "000001000100", "000001000100", "000001000011", "000001000010", "000001000010", "000001000001", "000001000000", "000001000000", "000000111111", "000000111110", "000000111110", "000000111101", "000000111101", "000000111100", "000000111011", "000000111011", "000000111010", "000000111001", "000000111001", "000000111000", "000000111000", "000000110111", "000000110111", "000000110110", "000000110101", "000000110101", "000000110100", "000000110100", "000000110011", "000000110011", "000000110010", "000000110010", "000000110001", "000000110001", "000000110000", "000000110000", "000000101111", "000000101111", "000000101110", "000000101110", "000000101101", "000000101101", "000000101100", "000000101100", "000000101011", "000000101011", "000000101010", "000000101010", "000000101001", "000000101001", "000000101001", "000000101000", "000000101000", "000000100111", "000000100111", "000000100110", "000000100110", "000000100110", "000000100101", "000000100101", "000000100100", "000000100100", "000000100100", "000000100011", "000000100011", "000000100011", "000000100010", "000000100010", "000000100001", "000000100001", "000000100001", "000000100000", "000000100000", "000000100000", "000000011111", "000000011111", "000000011111", "000000011110", "000000011110", "000000011110", "000000011110", "000000011101", "000000011101", "000000011101", "000000011100", "000000011100", "000000011100", "000000011100", "000000011011", "000000011011", "000000011011", "000000011011", "000000011010", "000000011010", "000000011010", "000000011010", "000000011001", "000000011001", "000000011001", "000000011001", "000000011001", "000000011000", "000000011000", "000000011000", "000000011000", "000000011000", "000000011000", "000000010111", "000000010111", "000000010111", "000000010111", "000000010111", "000000010111", "000000010110", "000000010110", "000000010110", "000000010110", "000000010110", "000000010110", "000000010110", "000000010110", "000000010110", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010100", "000000010100", "000000010100", "000000010100", "000000010100", "000000010100", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010101", "000000010110", "000000010110", "000000010110", "000000010110", "000000010110", "000000010110", "000000010110", "000000010110", "000000010111", "000000010111", "000000010111", "000000010111", "000000010111", "000000010111", "000000010111", "000000011000", "000000011000", "000000011000", "000000011000", "000000011000", "000000011001", "000000011001", "000000011001", "000000011001", "000000011001", "000000011010", "000000011010", "000000011010", "000000011010", "000000011010", "000000011011", "000000011011", "000000011011", "000000011011", "000000011100", "000000011100", "000000011100", "000000011101", "000000011101", "000000011101", "000000011101", "000000011110", "000000011110", "000000011110", "000000011111", "000000011111", "000000011111", "000000100000", "000000100000", "000000100000", "000000100001", "000000100001", "000000100001", "000000100010", "000000100010", "000000100010", "000000100011", "000000100011", "000000100011", "000000100100", "000000100100", "000000100101", "000000100101", "000000100101", "000000100110", "000000100110", "000000100111", "000000100111", "000000100111", "000000101000", "000000101000", "000000101001", "000000101001", "000000101010", "000000101010", "000000101011", "000000101011", "000000101011", "000000101100", "000000101100", "000000101101", "000000101101", "000000101110", "000000101110", "000000101111", "000000101111", "000000110000", "000000110000", "000000110001", "000000110001", "000000110010", "000000110010", "000000110011", "000000110100", "000000110100", "000000110101", "000000110101", "000000110110", "000000110110", "000000110111", "000000110111", "000000111000", "000000111001", "000000111001", "000000111010", "000000111010", "000000111011", "000000111100", "000000111100", "000000111101", "000000111101", "000000111110", "000000111111", "000000111111", "000001000000", "000001000001", "000001000001", "000001000010", "000001000011", "000001000011", "000001000100", "000001000101", "000001000101", "000001000110", "000001000111", "000001000111", "000001001000", "000001001001", "000001001001", "000001001010", "000001001011", "000001001100", "000001001100", "000001001101", "000001001110", "000001001110", "000001001111", "000001010000", "000001010001", "000001010001", "000001010010", "000001010011", "000001010100", "000001010101", "000001010101", "000001010110", "000001010111", "000001011000", "000001011000", "000001011001", "000001011010", "000001011011", "000001011100", "000001011100", "000001011101", "000001011110", "000001011111", "000001100000", "000001100001", "000001100010", "000001100010", "000001100011", "000001100100", "000001100101", "000001100110", "000001100111", "000001101000", "000001101000", "000001101001", "000001101010", "000001101011", "000001101100", "000001101101", "000001101110", "000001101111", "000001110000", "000001110001", "000001110010", "000001110010", "000001110011", "000001110100", "000001110101", "000001110110", "000001110111", "000001111000", "000001111001", "000001111010", "000001111011", "000001111100", "000001111101", "000001111110", "000001111111", "000010000000", "000010000001", "000010000010", "000010000011", "000010000100", "000010000101", "000010000110", "000010000111", "000010001000", "000010001001", "000010001010", "000010001011", "000010001100", "000010001101", "000010001110", "000010010000", "000010010001", "000010010010", "000010010011", "000010010100", "000010010101", "000010010110", "000010010111", "000010011000", "000010011001", "000010011010", "000010011100", "000010011101", "000010011110", "000010011111", "000010100000", "000010100001", "000010100010", "000010100011", "000010100101", "000010100110", "000010100111", "000010101000", "000010101001", "000010101010", "000010101100", "000010101101", "000010101110", "000010101111", "000010110000", "000010110010", "000010110011", "000010110100", "000010110101", "000010110110", "000010111000", "000010111001", "000010111010", "000010111011", "000010111101", "000010111110", "000010111111", "000011000000", "000011000010", "000011000011", "000011000100", "000011000101", "000011000111", "000011001000", "000011001001", "000011001010", "000011001100", "000011001101", "000011001110", "000011010000", "000011010001", "000011010010", "000011010100", "000011010101", "000011010110", "000011011000", "000011011001", "000011011010", "000011011100", "000011011101", "000011011110", "000011100000", "000011100001", "000011100010", "000011100100", "000011100101", "000011100110", "000011101000", "000011101001", "000011101011", "000011101100", "000011101101", "000011101111", "000011110000", "000011110010", "000011110011", "000011110100", "000011110110", "000011110111", "000011111001", "000011111010", "000011111100", "000011111101", "000011111110", "000100000000", "000100000001", "000100000011", "000100000100", "000100000110", "000100000111", "000100001001", "000100001010", "000100001100", "000100001101", "000100001111", "000100010000", "000100010010", "000100010011", "000100010101", "000100010110", "000100011000", "000100011001", "000100011011", "000100011100", "000100011110", "000100011111", "000100100001", "000100100010", "000100100100", "000100100110", "000100100111", "000100101001", "000100101010", "000100101100", "000100101101", "000100101111", "000100110001", "000100110010", "000100110100", "000100110101", "000100110111", "000100111001", "000100111010", "000100111100", "000100111101", "000100111111", "000101000001", "000101000010", "000101000100", "000101000110", "000101000111", "000101001001", "000101001011", "000101001100", "000101001110", "000101010000", "000101010001", "000101010011", "000101010101", "000101010110", "000101011000", "000101011010", "000101011011", "000101011101", "000101011111", "000101100000", "000101100010", "000101100100", "000101100110", "000101100111", "000101101001", "000101101011", "000101101100", "000101101110", "000101110000", "000101110010", "000101110011", "000101110101", "000101110111", "000101111001", "000101111010", "000101111100", "000101111110", "000110000000", "000110000001", "000110000011", "000110000101", "000110000111", "000110001001", "000110001010", "000110001100", "000110001110", "000110010000", "000110010010", "000110010011", "000110010101", "000110010111", "000110011001", "000110011011", "000110011101", "000110011110", "000110100000", "000110100010", "000110100100", "000110100110", "000110101000", "000110101010", "000110101011", "000110101101", "000110101111", "000110110001", "000110110011", "000110110101", "000110110111", "000110111001", "000110111011", "000110111100", "000110111110", "000111000000", "000111000010", "000111000100", "000111000110", "000111001000", "000111001010", "000111001100", "000111001110", "000111010000", "000111010010", "000111010100", "000111010110", "000111010111", "000111011001", "000111011011", "000111011101", "000111011111", "000111100001", "000111100011", "000111100101", "000111100111", "000111101001", "000111101011", "000111101101", "000111101111", "000111110001", "000111110011", "000111110101", "000111110111", "000111111001", "000111111011", "000111111101", "000111111111", "001000000001", "001000000011", "001000000101", "001000000111", "001000001010", "001000001100", "001000001110", "001000010000", "001000010010", "001000010100", "001000010110", "001000011000", "001000011010", "001000011100", "001000011110", "001000100000", "001000100010", "001000100100", "001000100111", "001000101001", "001000101011", "001000101101", "001000101111", "001000110001", "001000110011", "001000110101", "001000110111", "001000111010", "001000111100", "001000111110", "001001000000", "001001000010", "001001000100", "001001000110", "001001001001", "001001001011", "001001001101", "001001001111", "001001010001", "001001010011", "001001010110", "001001011000", "001001011010", "001001011100", "001001011110", "001001100000", "001001100011", "001001100101", "001001100111", "001001101001", "001001101011", "001001101110", "001001110000", "001001110010", "001001110100", "001001110110", "001001111001", "001001111011", "001001111101", "001001111111", "001010000010", "001010000100", "001010000110", "001010001000", "001010001011", "001010001101", "001010001111", "001010010001", "001010010100", "001010010110", "001010011000", "001010011010", "001010011101", "001010011111", "001010100001", "001010100100", "001010100110", "001010101000", "001010101011", "001010101101", "001010101111", "001010110001", "001010110100", "001010110110", "001010111000", "001010111011", "001010111101", "001010111111", "001011000010", "001011000100", "001011000110", "001011001001", "001011001011", "001011001101", "001011010000", "001011010010", "001011010100", "001011010111", "001011011001", "001011011011", "001011011110", "001011100000", "001011100011", "001011100101", "001011100111", "001011101010", "001011101100", "001011101111", "001011110001", "001011110011", "001011110110", "001011111000", "001011111011", "001011111101", "001011111111", "001100000010", "001100000100", "001100000111", "001100001001", "001100001011", "001100001110", "001100010000", "001100010011", "001100010101", "001100011000", "001100011010", "001100011100", "001100011111", "001100100001", "001100100100", "001100100110", "001100101001", "001100101011", "001100101110", "001100110000", "001100110011", "001100110101", "001100111000", "001100111010", "001100111101", "001100111111", "001101000010", "001101000100", "001101000111", "001101001001", "001101001011", "001101001110", "001101010001", "001101010011", "001101010110", "001101011000", "001101011011", "001101011101", "001101100000", "001101100010", "001101100101", "001101100111", "001101101010", "001101101100", "001101101111", "001101110001", "001101110100", "001101110110", "001101111001", "001101111100", "001101111110", "001110000001", "001110000011", "001110000110", "001110001000", "001110001011", "001110001101", "001110010000", "001110010011", "001110010101", "001110011000", "001110011010", "001110011101", "001110100000", "001110100010", "001110100101", "001110100111", "001110101010", "001110101101", "001110101111", "001110110010", "001110110100", "001110110111", "001110111010", "001110111100", "001110111111", "001111000001", "001111000100", "001111000111", "001111001001", "001111001100", "001111001111", "001111010001", "001111010100", "001111010111", "001111011001", "001111011100", "001111011111", "001111100001", "001111100100", "001111100111", "001111101001", "001111101100", "001111101111", "001111110001", "001111110100", "001111110111", "001111111001", "001111111100", "001111111111", "010000000001", "010000000100", "010000000111", "010000001001", "010000001100", "010000001111", "010000010001", "010000010100", "010000010111", "010000011010", "010000011100", "010000011111", "010000100010", "010000100100", "010000100111", "010000101010", "010000101101", "010000101111", "010000110010", "010000110101", "010000110111", "010000111010", "010000111101", "010001000000", "010001000010", "010001000101", "010001001000", "010001001011", "010001001101", "010001010000", "010001010011", "010001010110", "010001011000", "010001011011", "010001011110", "010001100001", "010001100011", "010001100110", "010001101001", "010001101100", "010001101111", "010001110001", "010001110100", "010001110111", "010001111010", "010001111100", "010001111111", "010010000010", "010010000101", "010010001000", "010010001010", "010010001101", "010010010000", "010010010011", "010010010110", "010010011000", "010010011011", "010010011110", "010010100001", "010010100100", "010010100110", "010010101001", "010010101100", "010010101111", "010010110010", "010010110101", "010010110111", "010010111010", "010010111101", "010011000000", "010011000011", "010011000110", "010011001000", "010011001011", "010011001110", "010011010001", "010011010100", "010011010111", "010011011010", "010011011100", "010011011111", "010011100010", "010011100101", "010011101000", "010011101011", "010011101110", "010011110000", "010011110011", "010011110110", "010011111001", "010011111100", "010011111111", "010100000010", "010100000101", "010100000111", "010100001010", "010100001101", "010100010000", "010100010011", "010100010110", "010100011001", "010100011100", "010100011111", "010100100001", "010100100100", "010100100111", "010100101010", "010100101101", "010100110000", "010100110011", "010100110110", "010100111001", "010100111100", "010100111111", "010101000001", "010101000100", "010101000111", "010101001010", "010101001101", "010101010000", "010101010011", "010101010110", "010101011001", "010101011100", "010101011111", "010101100010", "010101100101", "010101101000", "010101101010", "010101101101", "010101110000", "010101110011", "010101110110", "010101111001", "010101111100", "010101111111", "010110000010", "010110000101", "010110001000", "010110001011", "010110001110", "010110010001", "010110010100", "010110010111", "010110011010", "010110011101", "010110100000", "010110100011", "010110100110", "010110101001", "010110101100", "010110101110", "010110110001", "010110110100", "010110110111", "010110111010", "010110111101", "010111000000", "010111000011", "010111000110", "010111001001", "010111001100", "010111001111", "010111010010", "010111010101", "010111011000", "010111011011", "010111011110", "010111100001", "010111100100", "010111100111", "010111101010", "010111101101", "010111110000", "010111110011", "010111110110", "010111111001", "010111111100", "010111111111", "011000000010", "011000000101", "011000001000", "011000001011", "011000001110", "011000010001", "011000010100", "011000010111", "011000011010", "011000011101", "011000100000", "011000100011", "011000100110", "011000101010", "011000101101", "011000110000", "011000110011", "011000110110", "011000111001", "011000111100", "011000111111", "011001000010", "011001000101", "011001001000", "011001001011", "011001001110", "011001010001", "011001010100", "011001010111", "011001011010", "011001011101", "011001100000", "011001100011", "011001100110", "011001101001", "011001101100", "011001101111", "011001110010", "011001110101", "011001111001", "011001111100", "011001111111", "011010000010", "011010000101", "011010001000", "011010001011", "011010001110", "011010010001", "011010010100", "011010010111", "011010011010", "011010011101", "011010100000", "011010100011", "011010100110", "011010101001", "011010101101", "011010110000", "011010110011", "011010110110", "011010111001", "011010111100", "011010111111", "011011000010", "011011000101", "011011001000", "011011001011", "011011001110", "011011010001", "011011010100", "011011011000", "011011011011", "011011011110", "011011100001", "011011100100", "011011100111", "011011101010", "011011101101", "011011110000", "011011110011", "011011110110", "011011111001", "011011111101", "011100000000", "011100000011", "011100000110", "011100001001", "011100001100", "011100001111", "011100010010", "011100010101", "011100011000", "011100011011", "011100011110", "011100100010", "011100100101", "011100101000", "011100101011", "011100101110", "011100110001", "011100110100", "011100110111", "011100111010", "011100111101", "011101000001", "011101000100", "011101000111", "011101001010", "011101001101", "011101010000", "011101010011", "011101010110", "011101011001", "011101011100", "011101011111", "011101100011", "011101100110", "011101101001", "011101101100", "011101101111", "011101110010", "011101110101", "011101111000", "011101111011", "011101111111", "011110000010", "011110000101", "011110001000", "011110001011", "011110001110", "011110010001", "011110010100", "011110010111", "011110011010", "011110011110", "011110100001", "011110100100", "011110100111", "011110101010", "011110101101", "011110110000", "011110110011", "011110110110", "011110111010", "011110111101", "011111000000", "011111000011", "011111000110", "011111001001", "011111001100", "011111001111", "011111010010", "011111010110", "011111011001", "011111011100", "011111011111", "011111100010", "011111100101", "011111101000", "011111101011", "011111101110", "011111110010", "011111110101", "011111111000", "011111111011", "011111111110", "100000000001", "100000000100", "100000000111", "100000001010", "100000001101", "100000010001", "100000010100", "100000010111", "100000011010", "100000011101", "100000100000", "100000100011", "100000100110", "100000101001", "100000101101", "100000110000", "100000110011", "100000110110", "100000111001", "100000111100", "100000111111", "100001000010", "100001000101", "100001001001", "100001001100", "100001001111", "100001010010", "100001010101", "100001011000", "100001011011", "100001011110", "100001100001", "100001100101", "100001101000", "100001101011", "100001101110", "100001110001", "100001110100", "100001110111", "100001111010", "100001111101", "100010000000", "100010000100", "100010000111", "100010001010", "100010001101", "100010010000", "100010010011", "100010010110", "100010011001", "100010011100", "100010100000", "100010100011", "100010100110", "100010101001", "100010101100", "100010101111", "100010110010", "100010110101", "100010111000", "100010111011", "100010111110", "100011000010", "100011000101", "100011001000", "100011001011", "100011001110", "100011010001", "100011010100", "100011010111", "100011011010", "100011011101", "100011100001", "100011100100", "100011100111", "100011101010", "100011101101", "100011110000", "100011110011", "100011110110", "100011111001", "100011111100", "100011111111", "100100000010", "100100000110", "100100001001", "100100001100", "100100001111", "100100010010", "100100010101", "100100011000", "100100011011", "100100011110", "100100100001", "100100100100", "100100100111", "100100101011", "100100101110", "100100110001", "100100110100", "100100110111", "100100111010", "100100111101", "100101000000", "100101000011", "100101000110", "100101001001", "100101001100", "100101001111", "100101010010", "100101010110", "100101011001", "100101011100", "100101011111", "100101100010", "100101100101", "100101101000", "100101101011", "100101101110", "100101110001", "100101110100", "100101110111", "100101111010", "100101111101", "100110000000", "100110000011", "100110000110", "100110001010", "100110001101", "100110010000", "100110010011", "100110010110", "100110011001", "100110011100", "100110011111", "100110100010", "100110100101", "100110101000", "100110101011", "100110101110", "100110110001", "100110110100", "100110110111", "100110111010", "100110111101", "100111000000", "100111000011", "100111000110", "100111001001", "100111001100", "100111001111", "100111010010", "100111010101", "100111011001", "100111011100", "100111011111", "100111100010", "100111100101", "100111101000", "100111101011", "100111101110", "100111110001", "100111110100", "100111110111", "100111111010", "100111111101", "101000000000", "101000000011", "101000000110", "101000001001", "101000001100", "101000001111", "101000010010", "101000010101", "101000011000", "101000011011", "101000011110", "101000100001", "101000100100", "101000100111", "101000101010", "101000101101", "101000110000", "101000110011", "101000110110", "101000111001", "101000111100", "101000111111", "101001000010", "101001000101", "101001001000", "101001001011", "101001001110", "101001010001", "101001010011", "101001010110", "101001011001", "101001011100", "101001011111", "101001100010", "101001100101", "101001101000", "101001101011", "101001101110", "101001110001", "101001110100", "101001110111", "101001111010", "101001111101", "101010000000", "101010000011", "101010000110", "101010001001", "101010001100", "101010001111", "101010010010", "101010010101", "101010010111", "101010011010", "101010011101", "101010100000", "101010100011", "101010100110", "101010101001", "101010101100", "101010101111", "101010110010", "101010110101", "101010111000", "101010111011", "101010111110", "101011000000", "101011000011", "101011000110", "101011001001", "101011001100", "101011001111", "101011010010", "101011010101", "101011011000", "101011011011", "101011011110", "101011100000", "101011100011", "101011100110", "101011101001", "101011101100", "101011101111", "101011110010", "101011110101", "101011111000", "101011111010", "101011111101", "101100000000", "101100000011", "101100000110", "101100001001", "101100001100", "101100001111", "101100010001", "101100010100", "101100010111", "101100011010", "101100011101", "101100100000", "101100100011", "101100100101", "101100101000", "101100101011", "101100101110", "101100110001", "101100110100", "101100110111", "101100111001", "101100111100", "101100111111", "101101000010", "101101000101", "101101001000", "101101001010", "101101001101", "101101010000", "101101010011", "101101010110", "101101011001", "101101011011", "101101011110", "101101100001", "101101100100", "101101100111", "101101101001", "101101101100", "101101101111", "101101110010", "101101110101", "101101110111", "101101111010", "101101111101", "101110000000", "101110000011", "101110000101", "101110001000", "101110001011", "101110001110", "101110010000", "101110010011", "101110010110", "101110011001", "101110011100", "101110011110", "101110100001", "101110100100", "101110100111", "101110101001", "101110101100", "101110101111", "101110110010", "101110110100", "101110110111", "101110111010", "101110111101", "101110111111", "101111000010", "101111000101", "101111001000", "101111001010", "101111001101", "101111010000", "101111010010", "101111010101", "101111011000", "101111011011", "101111011101", "101111100000", "101111100011", "101111100101", "101111101000", "101111101011", "101111101110", "101111110000", "101111110011", "101111110110", "101111111000", "101111111011", "101111111110", "110000000000", "110000000011", "110000000110", "110000001000", "110000001011", "110000001110", "110000010000", "110000010011", "110000010110", "110000011000", "110000011011", "110000011110", "110000100000", "110000100011", "110000100110", "110000101000", "110000101011", "110000101110", "110000110000", "110000110011", "110000110110", "110000111000", "110000111011", "110000111110", "110001000000", "110001000011", "110001000101", "110001001000", "110001001011", "110001001101", "110001010000", "110001010010", "110001010101", "110001011000", "110001011010", "110001011101", "110001011111", "110001100010", "110001100101", "110001100111", "110001101010", "110001101100", "110001101111", "110001110010", "110001110100", "110001110111", "110001111001", "110001111100", "110001111110", "110010000001", "110010000011", "110010000110", "110010001001", "110010001011", "110010001110", "110010010000", "110010010011", "110010010101", "110010011000", "110010011010", "110010011101", "110010011111", "110010100010", "110010100100", "110010100111", "110010101001", "110010101100", "110010101110", "110010110001", "110010110100", "110010110110", "110010111000", "110010111011", "110010111101", "110011000000", "110011000010", "110011000101", "110011000111", "110011001010", "110011001100", "110011001111", "110011010001", "110011010100", "110011010110", "110011011001", "110011011011", "110011011110", "110011100000", "110011100011", "110011100101", "110011100111", "110011101010", "110011101100", "110011101111", "110011110001", "110011110100", "110011110110", "110011111000", "110011111011", "110011111101", "110100000000", "110100000010", "110100000100", "110100000111", "110100001001", "110100001100", "110100001110", "110100010000", "110100010011", "110100010101", "110100011000", "110100011010", "110100011100", "110100011111", "110100100001", "110100100100", "110100100110", "110100101000", "110100101011", "110100101101", "110100101111", "110100110010", "110100110100", "110100110110", "110100111001", "110100111011", "110100111101", "110101000000", "110101000010", "110101000100", "110101000111", "110101001001", "110101001011", "110101001110", "110101010000", "110101010010", "110101010100", "110101010111", "110101011001", "110101011011", "110101011110", "110101100000", "110101100010", "110101100101", "110101100111", "110101101001", "110101101011", "110101101110", "110101110000", "110101110010", "110101110100", "110101110111", "110101111001", "110101111011", "110101111101", "110110000000", "110110000010", "110110000100", "110110000110", "110110001001", "110110001011", "110110001101", "110110001111", "110110010001", "110110010100", "110110010110", "110110011000", "110110011010", "110110011100", "110110011111", "110110100001", "110110100011", "110110100101", "110110100111", "110110101001", "110110101100", "110110101110", "110110110000", "110110110010", "110110110100", "110110110110", "110110111001", "110110111011", "110110111101", "110110111111", "110111000001", "110111000011", "110111000101", "110111001000", "110111001010", "110111001100", "110111001110", "110111010000", "110111010010", "110111010100", "110111010110", "110111011000", "110111011011", "110111011101", "110111011111", "110111100001", "110111100011", "110111100101", "110111100111", "110111101001", "110111101011", "110111101101", "110111101111", "110111110001", "110111110011", "110111110101", "110111111000", "110111111010", "110111111100", "110111111110", "111000000000", "111000000010", "111000000100", "111000000110", "111000001000", "111000001010", "111000001100", "111000001110", "111000010000", "111000010010", "111000010100", "111000010110", "111000011000", "111000011010", "111000011100", "111000011110", "111000100000", "111000100010", "111000100100", "111000100110", "111000101000", "111000101001", "111000101011", "111000101101", "111000101111", "111000110001", "111000110011", "111000110101", "111000110111", "111000111001", "111000111011", "111000111101", "111000111111", "111001000001", "111001000011", "111001000100", "111001000110", "111001001000", "111001001010", "111001001100", "111001001110", "111001010000", "111001010010", "111001010100", "111001010101", "111001010111", "111001011001", "111001011011", "111001011101", "111001011111", "111001100001", "111001100010", "111001100100", "111001100110", "111001101000", "111001101010", "111001101100", "111001101101", "111001101111", "111001110001", "111001110011", "111001110101", "111001110110", "111001111000", "111001111010", "111001111100", "111001111110", "111001111111", "111010000001", "111010000011", "111010000101", "111010000110", "111010001000", "111010001010", "111010001100", "111010001101", "111010001111", "111010010001", "111010010011", "111010010100", "111010010110", "111010011000", "111010011001", "111010011011", "111010011101", "111010011111", "111010100000", "111010100010", "111010100100", "111010100101", "111010100111", "111010101001", "111010101010", "111010101100", "111010101110", "111010101111", "111010110001", "111010110011", "111010110100", "111010110110", "111010111000", "111010111001", "111010111011", "111010111101", "111010111110", "111011000000", "111011000010", "111011000011", "111011000101", "111011000110", "111011001000", "111011001010", "111011001011", "111011001101", "111011001110", "111011010000", "111011010010", "111011010011", "111011010101", "111011010110", "111011011000", "111011011001", "111011011011", "111011011101", "111011011110", "111011100000", "111011100001", "111011100011", "111011100100", "111011100110", "111011100111", "111011101001", "111011101010", "111011101100", "111011101101", "111011101111", "111011110000", "111011110010", "111011110011", "111011110101", "111011110110", "111011111000", "111011111001", "111011111011", "111011111100", "111011111110", "111011111111", "111100000001", "111100000010", "111100000011", "111100000101", "111100000110", "111100001000", "111100001001", "111100001011", "111100001100", "111100001101", "111100001111", "111100010000", "111100010010", "111100010011", "111100010100", "111100010110", "111100010111", "111100011001", "111100011010", "111100011011", "111100011101", "111100011110", "111100011111", "111100100001", "111100100010", "111100100011", "111100100101", "111100100110", "111100100111", "111100101001", "111100101010", "111100101011", "111100101101", "111100101110", "111100101111", "111100110001", "111100110010", "111100110011", "111100110101", "111100110110", "111100110111", "111100111000", "111100111010", "111100111011", "111100111100", "111100111101", "111100111111", "111101000000", "111101000001", "111101000010", "111101000100", "111101000101", "111101000110", "111101000111", "111101001001", "111101001010", "111101001011", "111101001100", "111101001101", "111101001111", "111101010000", "111101010001", "111101010010", "111101010011", "111101010101", "111101010110", "111101010111", "111101011000", "111101011001", "111101011010", "111101011100", "111101011101", "111101011110", "111101011111", "111101100000", "111101100001", "111101100010", "111101100011", "111101100101", "111101100110", "111101100111", "111101101000", "111101101001", "111101101010", "111101101011", "111101101100", "111101101101", "111101101110", "111101101111", "111101110001", "111101110010", "111101110011", "111101110100", "111101110101", "111101110110", "111101110111", "111101111000", "111101111001", "111101111010", "111101111011", "111101111100", "111101111101", "111101111110", "111101111111", "111110000000", "111110000001", "111110000010", "111110000011", "111110000100", "111110000101", "111110000110", "111110000111", "111110001000", "111110001001", "111110001010", "111110001011", "111110001100", "111110001101", "111110001101", "111110001110", "111110001111", "111110010000", "111110010001", "111110010010", "111110010011", "111110010100", "111110010101", "111110010110", "111110010111", "111110010111", "111110011000", "111110011001", "111110011010", "111110011011", "111110011100", "111110011101", "111110011101", "111110011110", "111110011111", "111110100000", "111110100001", "111110100010", "111110100011", "111110100011", "111110100100", "111110100101", "111110100110", "111110100111", "111110100111", "111110101000", "111110101001", "111110101010", "111110101010", "111110101011", "111110101100", "111110101101", "111110101110", "111110101110", "111110101111", "111110110000", "111110110001", "111110110001", "111110110010", "111110110011", "111110110011", "111110110100", "111110110101", "111110110110", "111110110110", "111110110111", "111110111000", "111110111000", "111110111001", "111110111010", "111110111010", "111110111011", "111110111100", "111110111100", "111110111101", "111110111110", "111110111110", "111110111111", "111111000000", "111111000000", "111111000001", "111111000010", "111111000010", "111111000011", "111111000011", "111111000100", "111111000101", "111111000101", "111111000110", "111111000110", "111111000111", "111111001000", "111111001000", "111111001001", "111111001001", "111111001010", "111111001010", "111111001011", "111111001011", "111111001100", "111111001101", "111111001101", "111111001110", "111111001110", "111111001111", "111111001111", "111111010000", "111111010000", "111111010001", "111111010001", "111111010010", "111111010010", "111111010011", "111111010011", "111111010100", "111111010100", "111111010100", "111111010101", "111111010101", "111111010110", "111111010110", "111111010111", "111111010111", "111111011000", "111111011000", "111111011000", "111111011001", "111111011001", "111111011010", "111111011010", "111111011010", "111111011011", "111111011011", "111111011100", "111111011100", "111111011100", "111111011101", "111111011101", "111111011101", "111111011110", "111111011110", "111111011110", "111111011111", "111111011111", "111111011111", "111111100000", "111111100000", "111111100000", "111111100001", "111111100001", "111111100001", "111111100010", "111111100010", "111111100010", "111111100010", "111111100011", "111111100011", "111111100011", "111111100100", "111111100100", "111111100100", "111111100100", "111111100101", "111111100101", "111111100101", "111111100101", "111111100101", "111111100110", "111111100110", "111111100110", "111111100110", "111111100110", "111111100111", "111111100111", "111111100111", "111111100111", "111111100111", "111111101000", "111111101000", "111111101000", "111111101000", "111111101000", "111111101000", "111111101000", "111111101001", "111111101001", "111111101001", "111111101001", "111111101001", "111111101001", "111111101001", "111111101001", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101011", "111111101011", "111111101011", "111111101011", "111111101011", "111111101011", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101010", "111111101001", "111111101001", "111111101001", "111111101001", "111111101001", "111111101001", "111111101001", "111111101001", "111111101001", "111111101000", "111111101000", "111111101000", "111111101000", "111111101000", "111111101000", "111111100111", "111111100111", "111111100111", "111111100111", "111111100111", "111111100111", "111111100110", "111111100110", "111111100110", "111111100110", "111111100110", "111111100101", "111111100101", "111111100101", "111111100101", "111111100100", "111111100100", "111111100100", "111111100100", "111111100011", "111111100011", "111111100011", "111111100011", "111111100010", "111111100010", "111111100010", "111111100001", "111111100001", "111111100001", "111111100001", "111111100000", "111111100000", "111111100000", "111111011111", "111111011111", "111111011111", "111111011110", "111111011110", "111111011110", "111111011101", "111111011101", "111111011100", "111111011100", "111111011100", "111111011011", "111111011011", "111111011011", "111111011010", "111111011010", "111111011001", "111111011001", "111111011001", "111111011000", "111111011000", "111111010111", "111111010111", "111111010110", "111111010110", "111111010110", "111111010101", "111111010101", "111111010100", "111111010100", "111111010011", "111111010011", "111111010010", "111111010010", "111111010001", "111111010001", "111111010000", "111111010000", "111111001111", "111111001111", "111111001110", "111111001110", "111111001101", "111111001101", "111111001100", "111111001100", "111111001011", "111111001011", "111111001010", "111111001010", "111111001001", "111111001000", "111111001000", "111111000111", "111111000111", "111111000110", "111111000110", "111111000101", "111111000100", "111111000100", "111111000011", "111111000010", "111111000010", "111111000001", "111111000001", "111111000000", "111110111111", "111110111111", "111110111110", "111110111101", "111110111101", "111110111100", "111110111011", "111110111011", "111110111010", "111110111001", "111110111001", "111110111000", "111110110111", "111110110111", "111110110110", "111110110101", "111110110101", "111110110100", "111110110011", "111110110010", "111110110010", "111110110001", "111110110000", "111110101111", "111110101111", "111110101110", "111110101101", "111110101100", "111110101100", "111110101011", "111110101010", "111110101001", "111110101001", "111110101000", "111110100111", "111110100110", "111110100101", "111110100101", "111110100100", "111110100011", "111110100010", "111110100001", "111110100000", "111110100000", "111110011111", "111110011110", "111110011101", "111110011100", "111110011011", "111110011010", "111110011010", "111110011001", "111110011000", "111110010111", "111110010110", "111110010101", "111110010100", "111110010011", "111110010011", "111110010010", "111110010001", "111110010000", "111110001111", "111110001110", "111110001101", "111110001100", "111110001011", "111110001010", "111110001001", "111110001000", "111110000111", "111110000110", "111110000101", "111110000100", "111110000011", "111110000010", "111110000001", "111110000000", "111101111111", "111101111110", "111101111101", "111101111100", "111101111011", "111101111010", "111101111001", "111101111000", "111101110111", "111101110110", "111101110101", "111101110100", "111101110011", "111101110010", "111101110001", "111101110000", "111101101111", "111101101110", "111101101101", "111101101100", "111101101011", "111101101010", "111101101000", "111101100111", "111101100110", "111101100101", "111101100100", "111101100011", "111101100010", "111101100001", "111101100000", "111101011110", "111101011101", "111101011100", "111101011011", "111101011010", "111101011001", "111101011000", "111101010110", "111101010101", "111101010100", "111101010011", "111101010010", "111101010000", "111101001111", "111101001110", "111101001101", "111101001100", "111101001010", "111101001001", "111101001000", "111101000111", "111101000110", "111101000100", "111101000011", "111101000010", "111101000001", "111100111111", "111100111110", "111100111101", "111100111100", "111100111010", "111100111001", "111100111000", "111100110111", "111100110101", "111100110100", "111100110011", "111100110001", "111100110000", "111100101111", "111100101101", "111100101100", "111100101011", "111100101001", "111100101000", "111100100111", "111100100101", "111100100100", "111100100011", "111100100001", "111100100000", "111100011111", "111100011101", "111100011100", "111100011011", "111100011001", "111100011000", "111100010111", "111100010101", "111100010100", "111100010010", "111100010001", "111100010000", "111100001110", "111100001101", "111100001011", "111100001010", "111100001000", "111100000111", "111100000110", "111100000100", "111100000011", "111100000001", "111100000000", "111011111110", "111011111101", "111011111011", "111011111010", "111011111000", "111011110111", "111011110110", "111011110100", "111011110011", "111011110001", "111011110000", "111011101110", "111011101101", "111011101011", "111011101010", "111011101000", "111011100111", "111011100101", "111011100011", "111011100010", "111011100000", "111011011111", "111011011101", "111011011100", "111011011010", "111011011001", "111011010111", "111011010101", "111011010100", "111011010010", "111011010001", "111011001111", "111011001110", "111011001100", "111011001010", "111011001001", "111011000111", "111011000110", "111011000100", "111011000010", "111011000001", "111010111111", "111010111101", "111010111100", "111010111010", "111010111001", "111010110111", "111010110101", "111010110100", "111010110010", "111010110000", "111010101111", "111010101101", "111010101011", "111010101010", "111010101000", "111010100110", "111010100101", "111010100011", "111010100001", "111010011111", "111010011110", "111010011100", "111010011010", "111010011001", "111010010111", "111010010101", "111010010011", "111010010010", "111010010000", "111010001110", "111010001100", "111010001011", "111010001001", "111010000111", "111010000101", "111010000100", "111010000010", "111010000000", "111001111110", "111001111101", "111001111011", "111001111001", "111001110111", "111001110101", "111001110100", "111001110010", "111001110000", "111001101110", "111001101100", "111001101011", "111001101001", "111001100111", "111001100101", "111001100011", "111001100001", "111001100000", "111001011110", "111001011100", "111001011010", "111001011000", "111001010110", "111001010100", "111001010011", "111001010001", "111001001111", "111001001101", "111001001011", "111001001001", "111001000111", "111001000101", "111001000011", "111001000010", "111001000000", "111000111110", "111000111100", "111000111010", "111000111000", "111000110110", "111000110100", "111000110010", "111000110000", "111000101110", "111000101100", "111000101010", "111000101001", "111000100111", "111000100101", "111000100011", "111000100001", "111000011111", "111000011101", "111000011011", "111000011001", "111000010111", "111000010101", "111000010011", "111000010001", "111000001111", "111000001101", "111000001011", "111000001001", "111000000111", "111000000101", "111000000011", "111000000001", "110111111111", "110111111101", "110111111011", "110111111001", "110111110111", "110111110100", "110111110010", "110111110000", "110111101110", "110111101100", "110111101010", "110111101000", "110111100110", "110111100100", "110111100010", "110111100000", "110111011110", "110111011100", "110111011010", "110111010111", "110111010101", "110111010011", "110111010001", "110111001111", "110111001101", "110111001011", "110111001001", "110111000111", "110111000100", "110111000010", "110111000000", "110110111110", "110110111100", "110110111010", "110110111000", "110110110101", "110110110011", "110110110001", "110110101111", "110110101101", "110110101011", "110110101000", "110110100110", "110110100100", "110110100010", "110110100000", "110110011101", "110110011011", "110110011001", "110110010111", "110110010101", "110110010010", "110110010000", "110110001110", "110110001100", "110110001010", "110110000111", "110110000101", "110110000011", "110110000001", "110101111110", "110101111100", "110101111010", "110101111000", "110101110101", "110101110011", "110101110001", "110101101111", "110101101100", "110101101010", "110101101000", "110101100110", "110101100011", "110101100001", "110101011111", "110101011101", "110101011010", "110101011000", "110101010110", "110101010011", "110101010001", "110101001111", "110101001100", "110101001010", "110101001000", "110101000101", "110101000011", "110101000001", "110100111111", "110100111100", "110100111010", "110100110111", "110100110101", "110100110011", "110100110000", "110100101110", "110100101100", "110100101001", "110100100111", "110100100101", "110100100010", "110100100000", "110100011110", "110100011011", "110100011001", "110100010110", "110100010100", "110100010010", "110100001111", "110100001101", "110100001010", "110100001000", "110100000110", "110100000011", "110100000001", "110011111110", "110011111100", "110011111010", "110011110111", "110011110101", "110011110010", "110011110000", "110011101110", "110011101011", "110011101001", "110011100110", "110011100100", "110011100001", "110011011111", "110011011100", "110011011010", "110011010111", "110011010101", "110011010011", "110011010000", "110011001110", "110011001011", "110011001001", "110011000110", "110011000100", "110011000001", "110010111111", "110010111100", "110010111010", "110010110111", "110010110101", "110010110010", "110010110000", "110010101101", "110010101011", "110010101000", "110010100110", "110010100011", "110010100001", "110010011110", "110010011100", "110010011001", "110010010111", "110010010100", "110010010001", "110010001111", "110010001100", "110010001010", "110010000111", "110010000101", "110010000010", "110010000000", "110001111101", "110001111010", "110001111000", "110001110101", "110001110011", "110001110000", "110001101110", "110001101011", "110001101000", "110001100110", "110001100011", "110001100001", "110001011110", "110001011100", "110001011001", "110001010110", "110001010100", "110001010001", "110001001111", "110001001100", "110001001001", "110001000111", "110001000100", "110001000001", "110000111111", "110000111100", "110000111010", "110000110111", "110000110100", "110000110010", "110000101111", "110000101100", "110000101010", "110000100111", "110000100100", "110000100010", "110000011111", "110000011100", "110000011010", "110000010111", "110000010100", "110000010010", "110000001111", "110000001100", "110000001010", "110000000111", "110000000100", "110000000010", "101111111111", "101111111100", "101111111010", "101111110111", "101111110100", "101111110010", "101111101111", "101111101100", "101111101010", "101111100111", "101111100100", "101111100001", "101111011111", "101111011100", "101111011001", "101111010111", "101111010100", "101111010001", "101111001110", "101111001100", "101111001001", "101111000110", "101111000011", "101111000001", "101110111110", "101110111011", "101110111001", "101110110110", "101110110011", "101110110000", "101110101110", "101110101011", "101110101000", "101110100101", "101110100010", "101110100000", "101110011101", "101110011010", "101110010111", "101110010101", "101110010010", "101110001111", "101110001100", "101110001010", "101110000111", "101110000100", "101110000001", "101101111110", "101101111100", "101101111001", "101101110110", "101101110011", "101101110000", "101101101110", "101101101011", "101101101000", "101101100101", "101101100010", "101101100000", "101101011101", "101101011010", "101101010111", "101101010100", "101101010001", "101101001111", "101101001100", "101101001001", "101101000110", "101101000011", "101101000000", "101100111110", "101100111011", "101100111000", "101100110101", "101100110010", "101100101111", "101100101101", "101100101010", "101100100111", "101100100100", "101100100001", "101100011110", "101100011011", "101100011001", "101100010110", "101100010011", "101100010000", "101100001101", "101100001010", "101100000111", "101100000101", "101100000010", "101011111111", "101011111100", "101011111001", "101011110110", "101011110011", "101011110000", "101011101101", "101011101011", "101011101000", "101011100101", "101011100010", "101011011111", "101011011100", "101011011001", "101011010110", "101011010011", "101011010000", "101011001110", "101011001011", "101011001000", "101011000101", "101011000010", "101010111111", "101010111100", "101010111001", "101010110110", "101010110011", "101010110000", "101010101101", "101010101011", "101010101000", "101010100101", "101010100010", "101010011111", "101010011100", "101010011001", "101010010110", "101010010011", "101010010000", "101010001101", "101010001010", "101010000111", "101010000100", "101010000001", "101001111110", "101001111011", "101001111001", "101001110110", "101001110011", "101001110000", "101001101101", "101001101010", "101001100111", "101001100100", "101001100001", "101001011110", "101001011011", "101001011000", "101001010101", "101001010010", "101001001111", "101001001100", "101001001001", "101001000110", "101001000011", "101001000000", "101000111101", "101000111010", "101000110111", "101000110100", "101000110001", "101000101110", "101000101011", "101000101000", "101000100101", "101000100010", "101000011111", "101000011100", "101000011001", "101000010110", "101000010011", "101000010000", "101000001101", "101000001010", "101000000111", "101000000100", "101000000001", "100111111110", "100111111011", "100111111000", "100111110101", "100111110010", "100111101111", "100111101100", "100111101001", "100111100110", "100111100011", "100111100000", "100111011101", "100111011010", "100111010111", "100111010100", "100111010001", "100111001110", "100111001011", "100111001000", "100111000101", "100111000010", "100110111111", "100110111100", "100110111001", "100110110110", "100110110011", "100110110000", "100110101101", "100110101010", "100110100110", "100110100011", "100110100000", "100110011101", "100110011010", "100110010111", "100110010100", "100110010001", "100110001110", "100110001011", "100110001000", "100110000101", "100110000010", "100101111111", "100101111100", "100101111001", "100101110110", "100101110011", "100101110000", "100101101100", "100101101001", "100101100110", "100101100011", "100101100000", "100101011101", "100101011010", "100101010111", "100101010100", "100101010001", "100101001110", "100101001011", "100101001000", "100101000101", "100101000010", "100100111111", "100100111011", "100100111000", "100100110101", "100100110010", "100100101111", "100100101100", "100100101001", "100100100110", "100100100011", "100100100000", "100100011101", "100100011010", "100100010111", "100100010011", "100100010000", "100100001101", "100100001010", "100100000111", "100100000100", "100100000001", "100011111110", "100011111011", "100011111000", "100011110101", "100011110010", "100011101110", "100011101011", "100011101000", "100011100101", "100011100010", "100011011111", "100011011100", "100011011001", "100011010110", "100011010011", "100011010000", "100011001100", "100011001001", "100011000110", "100011000011", "100011000000", "100010111101", "100010111010", "100010110111", "100010110100", "100010110001", "100010101101", "100010101010", "100010100111", "100010100100", "100010100001", "100010011110", "100010011011", "100010011000", "100010010101", "100010010010", "100010001110", "100010001011", "100010001000", "100010000101", "100010000010", "100001111111", "100001111100", "100001111001", "100001110110", "100001110011", "100001101111", "100001101100", "100001101001", "100001100110", "100001100011", "100001100000", "100001011101", "100001011010", "100001010111", "100001010011", "100001010000", "100001001101", "100001001010", "100001000111", "100001000100", "100001000001", "100000111110", "100000111011", "100000110111", "100000110100", "100000110001", "100000101110", "100000101011", "100000101000", "100000100101", "100000100010", "100000011111", "100000011011", "100000011000", "100000010101", "100000010010", "100000001111", "100000001100", "100000001001", "100000000110", "100000000011", "100000000000"
 );

signal counter_next : unsigned(11 downto 0) := (others => '0'); 
signal counter_sine_next : unsigned(11 downto 0) := (others => '0'); 
signal counter_reg : unsigned(11 downto 0) := (others => '0'); 
signal counter_sine_reg : unsigned(11 downto 0) := (others => '0'); 
signal sine_value_A, sine_value_B, sine_value_C : unsigned(11 downto 0) := (others => '0');  
signal gates : std_logic_vector(5 downto 0) := (others => '0'); 
signal igbt_in, igbt_out : std_logic_vector(5 downto 0) := (others => '0'); 
signal sine_tick, carrier_tick : std_logic;

begin
-- Componente divisor frecuencia contador modulo m
sine_modm_unit: entity work.modm(Behavioral)
    generic map(N => 16)
    port map(clk => clk, reset => reset, enable => enable_reg, q => open, max_tick => sine_tick, M => freq_sine);

carrier_modm_unit: entity work.modm(Behavioral)
    generic map(N => 16)
    port map(clk => clk, reset => reset, enable => enable_reg, q => open, max_tick => carrier_tick, M => freq_carrier);

delay_U_unit: entity work.retardo(Behavioral)
    port map(clk => clk, reset => reset, igbt_in => igbt_in(1 downto 0), igbt_out => igbt_out(1 downto 0));
    
delay_V_unit: entity work.retardo(Behavioral)
    port map(clk => clk, reset => reset, igbt_in => igbt_in(3 downto 2), igbt_out => igbt_out(3 downto 2));
    
delay_W_unit: entity work.retardo(Behavioral)
    port map(clk => clk, reset => reset, igbt_in => igbt_in(5 downto 4), igbt_out => igbt_out(5 downto 4));
    
       


-- register
process(clk, reset)
begin
    if reset = '1' then
        counter_reg <= (others => '0');
        counter_sine_reg <= (others => '0');
        enable_reg <= '0';
        state_reg <= '0';
    elsif rising_edge(clk) then
            counter_reg <= counter_next; 
            counter_sine_reg <= counter_sine_next; 
            enable_reg <= enable_next;
            state_reg <= state_next;
    end if;
end process;



process(start,state_reg,enable_reg, carrier_tick, sine_tick, counter_reg, counter_sine_reg)
begin
state_next <= state_reg;
counter_next <= counter_reg;
counter_sine_next <= counter_sine_reg;
enable_next <= enable_reg;
case state_reg is
    when '1' =>
        enable_next <= '1';
        if carrier_tick='1' then
            counter_next <= counter_reg+1;
        end if;
        if sine_tick='1' then
            counter_sine_next <= counter_sine_reg+1;
        end if;   
    when others =>
        enable_next <= '0';
        state_next <= '0';
        if start ='1' then
           enable_next <='1';
           state_next <= '1';
        end if;    
end case;
end process;

process(counter_reg, counter_sine_reg, sine_value_A, sine_value_B, sine_value_C)
begin
    sine_value_A <= sine_table(to_integer(unsigned(counter_sine_reg)));
    sine_value_B <= sine_table(to_integer(unsigned(counter_sine_reg + 1365))); -- Desfase de 120
    sine_value_C <= sine_table(to_integer(unsigned(counter_sine_reg + 2730))); -- Desfase de 240
    
    if counter_reg <  (sine_value_A) then
        gates(0) <= '1';
        gates(1) <= '0';
    else
        gates(0) <= '0';
        gates(1) <= '1';    
    end if;
    if counter_reg <  (sine_value_B) then
        gates(2) <= '1';
        gates(3) <= '0';
    else 
        gates(2) <= '0';
        gates(3) <= '1';    
    end if;
    if counter_reg <  (sine_value_C) then
        gates(4) <= '1';
        gates(5) <= '0';
    else
        gates(4) <= '0';
        gates(5) <= '1';    
    end if;
end process;

-- output logic
igbt_in <= gates when enable_reg='1' else "000000"; 
igbt <= igbt_out when mode='1' else "00" & igbt_out(1) & igbt_out(0) & igbt_out(0) & igbt_out(1);


LED(5 downto 0) <= igbt_out(5 downto 0); 
LED(13 downto 6) <=  (others => '0'); 
LED(15) <=  '1' when mode='1' else '0';
LED(14) <=  '1' when enable_reg='1' else '0';


enable <= enable_reg;

end Behavioral;
